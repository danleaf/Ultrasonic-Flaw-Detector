module packet();

endmodule
