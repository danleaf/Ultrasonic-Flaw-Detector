module gain
(
	input [7:0] i_data,
	output [7:0] o_da_data
);
	
	assign o_da_data = i_data;
	
endmodule
	